// Levi de Lima Pereira Júnior - 121210472
// Roteiro 5 

parameter divide_by=100000000;  // divisor do clock de referência
// A frequencia do clock de referencia é 50 MHz.
// A frequencia de clk_2 será de  50 MHz / divide_by

parameter NBITS_INSTR = 32;
parameter NBITS_TOP = 8, NREGS_TOP = 32, NBITS_LCD = 64;
module top(input  logic clk_2,
           input  logic [NBITS_TOP-1:0] SWI,
           output logic [NBITS_TOP-1:0] LED,
           output logic [NBITS_TOP-1:0] SEG,
           output logic [NBITS_LCD-1:0] lcd_a, lcd_b,
           output logic [NBITS_INSTR-1:0] lcd_instruction,
           output logic [NBITS_TOP-1:0] lcd_registrador [0:NREGS_TOP-1],
           output logic [NBITS_TOP-1:0] lcd_pc, lcd_SrcA, lcd_SrcB,
             lcd_ALUResult, lcd_Result, lcd_WriteData, lcd_ReadData, 
           output logic lcd_MemWrite, lcd_Branch, lcd_MemtoReg, lcd_RegWrite);

  always_comb begin
    lcd_WriteData <= SWI;
    lcd_pc <= 'h12;
    lcd_instruction <= 'h34567890;
    lcd_SrcA <= 'hab;
    lcd_SrcB <= 'hcd;
    lcd_ALUResult <= 'hef;
    lcd_Result <= 'h11;
    lcd_ReadData <= 'h33;
    lcd_MemWrite <= SWI[0];
    lcd_Branch <= SWI[1];
    lcd_MemtoReg <= SWI[2];
    lcd_RegWrite <= SWI[3];
    for(int i=0; i<NREGS_TOP; i++)
       if(i != NREGS_TOP/2-1) lcd_registrador[i] <= i+i*16;
       else                   lcd_registrador[i] <= ~SWI;
    lcd_a <= {56'h1234567890ABCD, SWI};
    lcd_b <= {SWI, 56'hFEDCBA09876543};
  end

  enum logic [3:0] {A, B, C, D} estado;
  logic [0:0] entradaSelecaoContagem;
  logic [7:4] entradaParalela;
  logic [0:0] entradaSerial;
  logic [0:0] bitSaida;
  logic [3:0] memoria;
  logic [0:0] reset;
  logic [0:0] load;

  always_comb entradaSelecaoContagem <= SWI[1];
  always_comb entradaParalela <= SWI[7:4];
  always_comb entradaSerial <= SWI[3];
  always_comb reset <= SWI[0];
  always_comb load <= SWI[2];
  
  always_ff @( posedge reset or posedge clk_2 ) begin
    if (reset) begin
        memoria <= 0;
    end else 
    if (load) begin
        memoria <= entradaParalela;
    end else 
    if (entradaSelecaoContagem) begin
        memoria <= memoria - 1;
    end
    else begin
        memoria <= memoria + 1;
    end

    case (memoria) 
        'b0000: SEG <= 'b00111111;
        'b0001: SEG <= 'b00000110;
        'b0010: SEG <= 'b01011011;
        'b0011: SEG <= 'b01001111;
        'b0100: SEG <= 'b01100110;
        'b0101: SEG <= 'b01101101;
        'b0110: SEG <= 'b01111101;
        'b0111: SEG <= 'b00000111;
        'b1000: SEG <= 'b01111111;
        'b1001: SEG <= 'b01100111;
        'b1010: SEG <= 'b01110111;
        'b1011: SEG <= 'b01111100;
        'b1100: SEG <= 'b00111001;
        'b1101: SEG <= 'b01011110;
        'b1110: SEG <= 'b01111001;
        'b1111: SEG <= 'b01110001;
    endcase
  end

  always_ff @(posedge clk_2) begin
    if (reset) begin
      estado <= A;
    end
    else begin
      unique case (estado)
        A:
          if (entradaSerial == 0) begin
            estado <= A;
          end
          else begin
            estado <= B;
          end
        B:
          if (entradaSerial == 0) begin
            estado <= A;
          end
          else begin
            estado <= C;
          end
        C:
          if (entradaSerial == 0) begin
            estado <= A;
          end
          else begin
            estado <= D;
          end
        D:
          if (entradaSerial == 0) begin
            estado <= A;
          end
          else begin
            estado <= D;
          end
      endcase
    end
  end

  always_comb bitSaida <= (estado == D);
  always_comb LED[0] <= bitSaida;
  always_comb LED[7] <= clk_2;
endmodule
